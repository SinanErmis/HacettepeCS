`timescale 1ns/10ps

module full_adder(
    input A, B, Cin,
    output S, Cout
);

	// Your code goes here.  DO NOT change anything that is already given! Otherwise, you will not be able to pass the tests!

endmodule
