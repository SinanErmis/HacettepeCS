`timescale 1 ns/10 ps

module four_bit_rca_tb;
	// Your code goes here.  DO NOT change anything that is already given! Otherwise, you will not be able to pass the tests!
endmodule