`timescale 1ns/10ps

module multiplier (
    input [2:0] A, B,
    output [5:0] P
);

	// Your code goes here.  DO NOT change anything that is already given! Otherwise, you will not be able to pass the tests!


endmodule
