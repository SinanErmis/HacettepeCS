module four_bit_rca(
    input [3:0] A,
    input [3:0] B,
    input Cin,
    output [3:0] S,
    output Cout
);
	// Your code goes here.  DO NOT change anything that is already given! Otherwise, you will not be able to pass the tests!
endmodule